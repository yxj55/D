module ysyx_25030093_addi(
    input clk,
    input rd_addr,
    input rs1_addr,
    input imm_data
    );
    wire 
    

endmodule