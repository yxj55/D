module ysyx_25030093_IFU(
    input [7:0] pc,
    input [31:0] inst
);
    ysyx_25030093_IDU u_ysyx_25030093_IDU(inst);
endmodule